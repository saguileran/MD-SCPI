<div id="toc_container">
  <p id="toc" class="toc_title" style="margin-top:-4px;">Table of Contents</p>
   <ul class="toc_list">
    <li><a href="#overview">Overview</a></li>
    <li><a href="#objectives">Objectives</a></li>
    <li><a href="#links-of-interest">Links of Interest</a></li>
    <li><a href="#weekly-reports">Weekly Reports</a></li>
    <li><a href="#output-files">Output Files</a></li>
    <li><a href="#references">References</a></li>
      <ul>
        <li><a href="#proteins-and-ligands">Proteins and Ligands</a></li>
        <li><a href="#software">Software</a></li>
      </ul>
    </ul>
</div>



<table rules="groups">
  <thead>
    <tr>
      <th style="text-align: left">Residue</th>
      <th style="text-align: center">Atom Numberth>
      <th style="text-align: right">AS4</th>
      <th style="text-align: right">COL</th>
    </tr>
  </thead>
  <tbody>
    <tr>
      <td style="text-align: left">SER</td>
      <td style="text-align: center">85</td>
      <td style="text-align: right">~</td>
      <td style="text-align: right"></td>
    </tr>
    <tr>
      <td style="text-align: left">ARGtd>
      <td style="text-align: center">92/td>
      <td style="text-align: right">*230</td>
      <td style="text-align: right"></td>
    </tr>
  </tbody>
  <tbody>
    <tr>
      <td style="text-align: left">GLN</td>
      <td style="text-align: center">51</td>
      <td style="text-align: right">*</td>
      <td style="text-align: right"></td>
    </tr>
    <tr>
      <td style="text-align: left">ASN</td>
      <td style="text-align: center">45</td>
      <td style="text-align: right"></td>
      <td style="text-align: right"></td>
    </tr>
  </tbody>
  <tbody>
    <tr>
      <td style="text-align: left">THR</td>
      <td style="text-align: center">220</td>
      <td style="text-align: right"></td>
      <td style="text-align: right"></td>
    </tr>
    <tr>
      <td style="text-align: left">HH</td>
      <td style="text-align: center">22</td>
      <td style="text-align: right"></td>
      <td style="text-align: right"></td>
    </tr>
  </tbody>
  <tbody>
    <tr>
      <td style="text-align: left">SER</td>
      <td style="text-align: center">118</td>
      <td style="text-align: right"></td>
      <td style="text-align: right"></td>
    </tr>
  </tbody>
<!--
  <tfoot>
    <tr>
      <td style="text-align: left">SER</td>
      <td style="text-align: center">118</td>
      <td style="text-align: right"></td>
      <td style="text-align: right"></td>
    </tr>
  </tfoot>
-->
</table>
  

